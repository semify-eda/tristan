package custom_instr_pkg;

  typedef enum logic [6:0] {
                            OPCODE_CNTB = 7'h6b,
                            OPCODE_WBITS = 7'h07
                            } cust_opcodes_e;

endpackage
  
